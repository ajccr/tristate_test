magic
tech sky130A
magscale 1 2
timestamp 1729812447
<< checkpaint >>
rect -3932 2548 23932 17660
<< viali >>
rect 6377 10625 6411 10659
rect 6561 10421 6595 10455
rect 6745 10081 6779 10115
rect 6377 10013 6411 10047
rect 6929 9945 6963 9979
rect 8585 9945 8619 9979
rect 6561 9877 6595 9911
rect 7481 9673 7515 9707
rect 7389 9537 7423 9571
<< metal1 >>
rect 6072 13626 13984 13648
rect 6072 13574 6886 13626
rect 6938 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 12886 13626
rect 12938 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 13984 13626
rect 6072 13552 13984 13574
rect 6072 13082 14012 13104
rect 6072 13030 7626 13082
rect 7678 13030 7690 13082
rect 7742 13030 7754 13082
rect 7806 13030 7818 13082
rect 7870 13030 7882 13082
rect 7934 13030 7946 13082
rect 7998 13030 13626 13082
rect 13678 13030 13690 13082
rect 13742 13030 13754 13082
rect 13806 13030 13818 13082
rect 13870 13030 13882 13082
rect 13934 13030 13946 13082
rect 13998 13030 14012 13082
rect 6072 13008 14012 13030
rect 6072 12538 13984 12560
rect 6072 12486 6886 12538
rect 6938 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 12886 12538
rect 12938 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 13984 12538
rect 6072 12464 13984 12486
rect 6072 11994 14012 12016
rect 6072 11942 7626 11994
rect 7678 11942 7690 11994
rect 7742 11942 7754 11994
rect 7806 11942 7818 11994
rect 7870 11942 7882 11994
rect 7934 11942 7946 11994
rect 7998 11942 13626 11994
rect 13678 11942 13690 11994
rect 13742 11942 13754 11994
rect 13806 11942 13818 11994
rect 13870 11942 13882 11994
rect 13934 11942 13946 11994
rect 13998 11942 14012 11994
rect 6072 11920 14012 11942
rect 6072 11450 13984 11472
rect 6072 11398 6886 11450
rect 6938 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 12886 11450
rect 12938 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 13984 11450
rect 6072 11376 13984 11398
rect 6072 10906 14012 10928
rect 6072 10854 7626 10906
rect 7678 10854 7690 10906
rect 7742 10854 7754 10906
rect 7806 10854 7818 10906
rect 7870 10854 7882 10906
rect 7934 10854 7946 10906
rect 7998 10854 13626 10906
rect 13678 10854 13690 10906
rect 13742 10854 13754 10906
rect 13806 10854 13818 10906
rect 13870 10854 13882 10906
rect 13934 10854 13946 10906
rect 13998 10854 14012 10906
rect 6072 10832 14012 10854
rect 6362 10616 6368 10668
rect 6420 10616 6426 10668
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6730 10452 6736 10464
rect 6595 10424 6736 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 6072 10362 13984 10384
rect 6072 10310 6886 10362
rect 6938 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 12886 10362
rect 12938 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 13984 10362
rect 6072 10288 13984 10310
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 4798 10004 4804 10056
rect 4856 10044 4862 10056
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 4856 10016 6377 10044
rect 4856 10004 4862 10016
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 6917 9979 6975 9985
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 7466 9976 7472 9988
rect 6963 9948 7472 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 8573 9979 8631 9985
rect 8573 9945 8585 9979
rect 8619 9976 8631 9979
rect 15194 9976 15200 9988
rect 8619 9948 15200 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 6549 9911 6607 9917
rect 6549 9877 6561 9911
rect 6595 9908 6607 9911
rect 7374 9908 7380 9920
rect 6595 9880 7380 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 6072 9818 14012 9840
rect 6072 9766 7626 9818
rect 7678 9766 7690 9818
rect 7742 9766 7754 9818
rect 7806 9766 7818 9818
rect 7870 9766 7882 9818
rect 7934 9766 7946 9818
rect 7998 9766 13626 9818
rect 13678 9766 13690 9818
rect 13742 9766 13754 9818
rect 13806 9766 13818 9818
rect 13870 9766 13882 9818
rect 13934 9766 13946 9818
rect 13998 9766 14012 9818
rect 6072 9744 14012 9766
rect 7466 9664 7472 9716
rect 7524 9664 7530 9716
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 6072 9274 13984 9296
rect 6072 9222 6886 9274
rect 6938 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 12886 9274
rect 12938 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 13984 9274
rect 6072 9200 13984 9222
rect 6072 8730 14012 8752
rect 6072 8678 7626 8730
rect 7678 8678 7690 8730
rect 7742 8678 7754 8730
rect 7806 8678 7818 8730
rect 7870 8678 7882 8730
rect 7934 8678 7946 8730
rect 7998 8678 13626 8730
rect 13678 8678 13690 8730
rect 13742 8678 13754 8730
rect 13806 8678 13818 8730
rect 13870 8678 13882 8730
rect 13934 8678 13946 8730
rect 13998 8678 14012 8730
rect 6072 8656 14012 8678
rect 6072 8186 13984 8208
rect 6072 8134 6886 8186
rect 6938 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 12886 8186
rect 12938 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 13984 8186
rect 6072 8112 13984 8134
rect 6072 7642 14012 7664
rect 6072 7590 7626 7642
rect 7678 7590 7690 7642
rect 7742 7590 7754 7642
rect 7806 7590 7818 7642
rect 7870 7590 7882 7642
rect 7934 7590 7946 7642
rect 7998 7590 13626 7642
rect 13678 7590 13690 7642
rect 13742 7590 13754 7642
rect 13806 7590 13818 7642
rect 13870 7590 13882 7642
rect 13934 7590 13946 7642
rect 13998 7590 14012 7642
rect 6072 7568 14012 7590
rect 6072 7098 13984 7120
rect 6072 7046 6886 7098
rect 6938 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 12886 7098
rect 12938 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 13984 7098
rect 6072 7024 13984 7046
rect 6072 6554 14012 6576
rect 6072 6502 7626 6554
rect 7678 6502 7690 6554
rect 7742 6502 7754 6554
rect 7806 6502 7818 6554
rect 7870 6502 7882 6554
rect 7934 6502 7946 6554
rect 7998 6502 13626 6554
rect 13678 6502 13690 6554
rect 13742 6502 13754 6554
rect 13806 6502 13818 6554
rect 13870 6502 13882 6554
rect 13934 6502 13946 6554
rect 13998 6502 14012 6554
rect 6072 6480 14012 6502
<< via1 >>
rect 6886 13574 6938 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 12886 13574 12938 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 7626 13030 7678 13082
rect 7690 13030 7742 13082
rect 7754 13030 7806 13082
rect 7818 13030 7870 13082
rect 7882 13030 7934 13082
rect 7946 13030 7998 13082
rect 13626 13030 13678 13082
rect 13690 13030 13742 13082
rect 13754 13030 13806 13082
rect 13818 13030 13870 13082
rect 13882 13030 13934 13082
rect 13946 13030 13998 13082
rect 6886 12486 6938 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 12886 12486 12938 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 7626 11942 7678 11994
rect 7690 11942 7742 11994
rect 7754 11942 7806 11994
rect 7818 11942 7870 11994
rect 7882 11942 7934 11994
rect 7946 11942 7998 11994
rect 13626 11942 13678 11994
rect 13690 11942 13742 11994
rect 13754 11942 13806 11994
rect 13818 11942 13870 11994
rect 13882 11942 13934 11994
rect 13946 11942 13998 11994
rect 6886 11398 6938 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 12886 11398 12938 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 7626 10854 7678 10906
rect 7690 10854 7742 10906
rect 7754 10854 7806 10906
rect 7818 10854 7870 10906
rect 7882 10854 7934 10906
rect 7946 10854 7998 10906
rect 13626 10854 13678 10906
rect 13690 10854 13742 10906
rect 13754 10854 13806 10906
rect 13818 10854 13870 10906
rect 13882 10854 13934 10906
rect 13946 10854 13998 10906
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 6736 10412 6788 10464
rect 6886 10310 6938 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 12886 10310 12938 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 4804 10004 4856 10056
rect 7472 9936 7524 9988
rect 15200 9936 15252 9988
rect 7380 9868 7432 9920
rect 7626 9766 7678 9818
rect 7690 9766 7742 9818
rect 7754 9766 7806 9818
rect 7818 9766 7870 9818
rect 7882 9766 7934 9818
rect 7946 9766 7998 9818
rect 13626 9766 13678 9818
rect 13690 9766 13742 9818
rect 13754 9766 13806 9818
rect 13818 9766 13870 9818
rect 13882 9766 13934 9818
rect 13946 9766 13998 9818
rect 7472 9707 7524 9716
rect 7472 9673 7481 9707
rect 7481 9673 7515 9707
rect 7515 9673 7524 9707
rect 7472 9664 7524 9673
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 6886 9222 6938 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 12886 9222 12938 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 7626 8678 7678 8730
rect 7690 8678 7742 8730
rect 7754 8678 7806 8730
rect 7818 8678 7870 8730
rect 7882 8678 7934 8730
rect 7946 8678 7998 8730
rect 13626 8678 13678 8730
rect 13690 8678 13742 8730
rect 13754 8678 13806 8730
rect 13818 8678 13870 8730
rect 13882 8678 13934 8730
rect 13946 8678 13998 8730
rect 6886 8134 6938 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 12886 8134 12938 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 7626 7590 7678 7642
rect 7690 7590 7742 7642
rect 7754 7590 7806 7642
rect 7818 7590 7870 7642
rect 7882 7590 7934 7642
rect 7946 7590 7998 7642
rect 13626 7590 13678 7642
rect 13690 7590 13742 7642
rect 13754 7590 13806 7642
rect 13818 7590 13870 7642
rect 13882 7590 13934 7642
rect 13946 7590 13998 7642
rect 6886 7046 6938 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 12886 7046 12938 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 7626 6502 7678 6554
rect 7690 6502 7742 6554
rect 7754 6502 7806 6554
rect 7818 6502 7870 6554
rect 7882 6502 7934 6554
rect 7946 6502 7998 6554
rect 13626 6502 13678 6554
rect 13690 6502 13742 6554
rect 13754 6502 13806 6554
rect 13818 6502 13870 6554
rect 13882 6502 13934 6554
rect 13946 6502 13998 6554
<< metal2 >>
rect 6884 13628 7260 13637
rect 6940 13626 6964 13628
rect 7020 13626 7044 13628
rect 7100 13626 7124 13628
rect 7180 13626 7204 13628
rect 6940 13574 6950 13626
rect 7194 13574 7204 13626
rect 6940 13572 6964 13574
rect 7020 13572 7044 13574
rect 7100 13572 7124 13574
rect 7180 13572 7204 13574
rect 6884 13563 7260 13572
rect 12884 13628 13260 13637
rect 12940 13626 12964 13628
rect 13020 13626 13044 13628
rect 13100 13626 13124 13628
rect 13180 13626 13204 13628
rect 12940 13574 12950 13626
rect 13194 13574 13204 13626
rect 12940 13572 12964 13574
rect 13020 13572 13044 13574
rect 13100 13572 13124 13574
rect 13180 13572 13204 13574
rect 12884 13563 13260 13572
rect 7624 13084 8000 13093
rect 7680 13082 7704 13084
rect 7760 13082 7784 13084
rect 7840 13082 7864 13084
rect 7920 13082 7944 13084
rect 7680 13030 7690 13082
rect 7934 13030 7944 13082
rect 7680 13028 7704 13030
rect 7760 13028 7784 13030
rect 7840 13028 7864 13030
rect 7920 13028 7944 13030
rect 7624 13019 8000 13028
rect 13624 13084 14000 13093
rect 13680 13082 13704 13084
rect 13760 13082 13784 13084
rect 13840 13082 13864 13084
rect 13920 13082 13944 13084
rect 13680 13030 13690 13082
rect 13934 13030 13944 13082
rect 13680 13028 13704 13030
rect 13760 13028 13784 13030
rect 13840 13028 13864 13030
rect 13920 13028 13944 13030
rect 13624 13019 14000 13028
rect 6884 12540 7260 12549
rect 6940 12538 6964 12540
rect 7020 12538 7044 12540
rect 7100 12538 7124 12540
rect 7180 12538 7204 12540
rect 6940 12486 6950 12538
rect 7194 12486 7204 12538
rect 6940 12484 6964 12486
rect 7020 12484 7044 12486
rect 7100 12484 7124 12486
rect 7180 12484 7204 12486
rect 6884 12475 7260 12484
rect 12884 12540 13260 12549
rect 12940 12538 12964 12540
rect 13020 12538 13044 12540
rect 13100 12538 13124 12540
rect 13180 12538 13204 12540
rect 12940 12486 12950 12538
rect 13194 12486 13204 12538
rect 12940 12484 12964 12486
rect 13020 12484 13044 12486
rect 13100 12484 13124 12486
rect 13180 12484 13204 12486
rect 12884 12475 13260 12484
rect 7624 11996 8000 12005
rect 7680 11994 7704 11996
rect 7760 11994 7784 11996
rect 7840 11994 7864 11996
rect 7920 11994 7944 11996
rect 7680 11942 7690 11994
rect 7934 11942 7944 11994
rect 7680 11940 7704 11942
rect 7760 11940 7784 11942
rect 7840 11940 7864 11942
rect 7920 11940 7944 11942
rect 7624 11931 8000 11940
rect 13624 11996 14000 12005
rect 13680 11994 13704 11996
rect 13760 11994 13784 11996
rect 13840 11994 13864 11996
rect 13920 11994 13944 11996
rect 13680 11942 13690 11994
rect 13934 11942 13944 11994
rect 13680 11940 13704 11942
rect 13760 11940 13784 11942
rect 13840 11940 13864 11942
rect 13920 11940 13944 11942
rect 13624 11931 14000 11940
rect 6884 11452 7260 11461
rect 6940 11450 6964 11452
rect 7020 11450 7044 11452
rect 7100 11450 7124 11452
rect 7180 11450 7204 11452
rect 6940 11398 6950 11450
rect 7194 11398 7204 11450
rect 6940 11396 6964 11398
rect 7020 11396 7044 11398
rect 7100 11396 7124 11398
rect 7180 11396 7204 11398
rect 6884 11387 7260 11396
rect 12884 11452 13260 11461
rect 12940 11450 12964 11452
rect 13020 11450 13044 11452
rect 13100 11450 13124 11452
rect 13180 11450 13204 11452
rect 12940 11398 12950 11450
rect 13194 11398 13204 11450
rect 12940 11396 12964 11398
rect 13020 11396 13044 11398
rect 13100 11396 13124 11398
rect 13180 11396 13204 11398
rect 12884 11387 13260 11396
rect 7624 10908 8000 10917
rect 7680 10906 7704 10908
rect 7760 10906 7784 10908
rect 7840 10906 7864 10908
rect 7920 10906 7944 10908
rect 7680 10854 7690 10906
rect 7934 10854 7944 10906
rect 7680 10852 7704 10854
rect 7760 10852 7784 10854
rect 7840 10852 7864 10854
rect 7920 10852 7944 10854
rect 7624 10843 8000 10852
rect 13624 10908 14000 10917
rect 13680 10906 13704 10908
rect 13760 10906 13784 10908
rect 13840 10906 13864 10908
rect 13920 10906 13944 10908
rect 13680 10854 13690 10906
rect 13934 10854 13944 10906
rect 13680 10852 13704 10854
rect 13760 10852 13784 10854
rect 13840 10852 13864 10854
rect 13920 10852 13944 10854
rect 13624 10843 14000 10852
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6380 10305 6408 10610
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6366 10296 6422 10305
rect 6366 10231 6422 10240
rect 6748 10130 6776 10406
rect 6884 10364 7260 10373
rect 6940 10362 6964 10364
rect 7020 10362 7044 10364
rect 7100 10362 7124 10364
rect 7180 10362 7204 10364
rect 6940 10310 6950 10362
rect 7194 10310 7204 10362
rect 6940 10308 6964 10310
rect 7020 10308 7044 10310
rect 7100 10308 7124 10310
rect 7180 10308 7204 10310
rect 6884 10299 7260 10308
rect 12884 10364 13260 10373
rect 12940 10362 12964 10364
rect 13020 10362 13044 10364
rect 13100 10362 13124 10364
rect 13180 10362 13204 10364
rect 12940 10310 12950 10362
rect 13194 10310 13204 10362
rect 12940 10308 12964 10310
rect 13020 10308 13044 10310
rect 13100 10308 13124 10310
rect 13180 10308 13204 10310
rect 12884 10299 13260 10308
rect 15198 10296 15254 10305
rect 15198 10231 15254 10240
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4816 9625 4844 9998
rect 15212 9994 15240 10231
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 4802 9616 4858 9625
rect 7392 9586 7420 9862
rect 7484 9722 7512 9930
rect 7624 9820 8000 9829
rect 7680 9818 7704 9820
rect 7760 9818 7784 9820
rect 7840 9818 7864 9820
rect 7920 9818 7944 9820
rect 7680 9766 7690 9818
rect 7934 9766 7944 9818
rect 7680 9764 7704 9766
rect 7760 9764 7784 9766
rect 7840 9764 7864 9766
rect 7920 9764 7944 9766
rect 7624 9755 8000 9764
rect 13624 9820 14000 9829
rect 13680 9818 13704 9820
rect 13760 9818 13784 9820
rect 13840 9818 13864 9820
rect 13920 9818 13944 9820
rect 13680 9766 13690 9818
rect 13934 9766 13944 9818
rect 13680 9764 13704 9766
rect 13760 9764 13784 9766
rect 13840 9764 13864 9766
rect 13920 9764 13944 9766
rect 13624 9755 14000 9764
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 4802 9551 4858 9560
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 6884 9276 7260 9285
rect 6940 9274 6964 9276
rect 7020 9274 7044 9276
rect 7100 9274 7124 9276
rect 7180 9274 7204 9276
rect 6940 9222 6950 9274
rect 7194 9222 7204 9274
rect 6940 9220 6964 9222
rect 7020 9220 7044 9222
rect 7100 9220 7124 9222
rect 7180 9220 7204 9222
rect 6884 9211 7260 9220
rect 12884 9276 13260 9285
rect 12940 9274 12964 9276
rect 13020 9274 13044 9276
rect 13100 9274 13124 9276
rect 13180 9274 13204 9276
rect 12940 9222 12950 9274
rect 13194 9222 13204 9274
rect 12940 9220 12964 9222
rect 13020 9220 13044 9222
rect 13100 9220 13124 9222
rect 13180 9220 13204 9222
rect 12884 9211 13260 9220
rect 7624 8732 8000 8741
rect 7680 8730 7704 8732
rect 7760 8730 7784 8732
rect 7840 8730 7864 8732
rect 7920 8730 7944 8732
rect 7680 8678 7690 8730
rect 7934 8678 7944 8730
rect 7680 8676 7704 8678
rect 7760 8676 7784 8678
rect 7840 8676 7864 8678
rect 7920 8676 7944 8678
rect 7624 8667 8000 8676
rect 13624 8732 14000 8741
rect 13680 8730 13704 8732
rect 13760 8730 13784 8732
rect 13840 8730 13864 8732
rect 13920 8730 13944 8732
rect 13680 8678 13690 8730
rect 13934 8678 13944 8730
rect 13680 8676 13704 8678
rect 13760 8676 13784 8678
rect 13840 8676 13864 8678
rect 13920 8676 13944 8678
rect 13624 8667 14000 8676
rect 6884 8188 7260 8197
rect 6940 8186 6964 8188
rect 7020 8186 7044 8188
rect 7100 8186 7124 8188
rect 7180 8186 7204 8188
rect 6940 8134 6950 8186
rect 7194 8134 7204 8186
rect 6940 8132 6964 8134
rect 7020 8132 7044 8134
rect 7100 8132 7124 8134
rect 7180 8132 7204 8134
rect 6884 8123 7260 8132
rect 12884 8188 13260 8197
rect 12940 8186 12964 8188
rect 13020 8186 13044 8188
rect 13100 8186 13124 8188
rect 13180 8186 13204 8188
rect 12940 8134 12950 8186
rect 13194 8134 13204 8186
rect 12940 8132 12964 8134
rect 13020 8132 13044 8134
rect 13100 8132 13124 8134
rect 13180 8132 13204 8134
rect 12884 8123 13260 8132
rect 7624 7644 8000 7653
rect 7680 7642 7704 7644
rect 7760 7642 7784 7644
rect 7840 7642 7864 7644
rect 7920 7642 7944 7644
rect 7680 7590 7690 7642
rect 7934 7590 7944 7642
rect 7680 7588 7704 7590
rect 7760 7588 7784 7590
rect 7840 7588 7864 7590
rect 7920 7588 7944 7590
rect 7624 7579 8000 7588
rect 13624 7644 14000 7653
rect 13680 7642 13704 7644
rect 13760 7642 13784 7644
rect 13840 7642 13864 7644
rect 13920 7642 13944 7644
rect 13680 7590 13690 7642
rect 13934 7590 13944 7642
rect 13680 7588 13704 7590
rect 13760 7588 13784 7590
rect 13840 7588 13864 7590
rect 13920 7588 13944 7590
rect 13624 7579 14000 7588
rect 6884 7100 7260 7109
rect 6940 7098 6964 7100
rect 7020 7098 7044 7100
rect 7100 7098 7124 7100
rect 7180 7098 7204 7100
rect 6940 7046 6950 7098
rect 7194 7046 7204 7098
rect 6940 7044 6964 7046
rect 7020 7044 7044 7046
rect 7100 7044 7124 7046
rect 7180 7044 7204 7046
rect 6884 7035 7260 7044
rect 12884 7100 13260 7109
rect 12940 7098 12964 7100
rect 13020 7098 13044 7100
rect 13100 7098 13124 7100
rect 13180 7098 13204 7100
rect 12940 7046 12950 7098
rect 13194 7046 13204 7098
rect 12940 7044 12964 7046
rect 13020 7044 13044 7046
rect 13100 7044 13124 7046
rect 13180 7044 13204 7046
rect 12884 7035 13260 7044
rect 7624 6556 8000 6565
rect 7680 6554 7704 6556
rect 7760 6554 7784 6556
rect 7840 6554 7864 6556
rect 7920 6554 7944 6556
rect 7680 6502 7690 6554
rect 7934 6502 7944 6554
rect 7680 6500 7704 6502
rect 7760 6500 7784 6502
rect 7840 6500 7864 6502
rect 7920 6500 7944 6502
rect 7624 6491 8000 6500
rect 13624 6556 14000 6565
rect 13680 6554 13704 6556
rect 13760 6554 13784 6556
rect 13840 6554 13864 6556
rect 13920 6554 13944 6556
rect 13680 6502 13690 6554
rect 13934 6502 13944 6554
rect 13680 6500 13704 6502
rect 13760 6500 13784 6502
rect 13840 6500 13864 6502
rect 13920 6500 13944 6502
rect 13624 6491 14000 6500
<< via2 >>
rect 6884 13626 6940 13628
rect 6964 13626 7020 13628
rect 7044 13626 7100 13628
rect 7124 13626 7180 13628
rect 7204 13626 7260 13628
rect 6884 13574 6886 13626
rect 6886 13574 6938 13626
rect 6938 13574 6940 13626
rect 6964 13574 7002 13626
rect 7002 13574 7014 13626
rect 7014 13574 7020 13626
rect 7044 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7100 13626
rect 7124 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7180 13626
rect 7204 13574 7206 13626
rect 7206 13574 7258 13626
rect 7258 13574 7260 13626
rect 6884 13572 6940 13574
rect 6964 13572 7020 13574
rect 7044 13572 7100 13574
rect 7124 13572 7180 13574
rect 7204 13572 7260 13574
rect 12884 13626 12940 13628
rect 12964 13626 13020 13628
rect 13044 13626 13100 13628
rect 13124 13626 13180 13628
rect 13204 13626 13260 13628
rect 12884 13574 12886 13626
rect 12886 13574 12938 13626
rect 12938 13574 12940 13626
rect 12964 13574 13002 13626
rect 13002 13574 13014 13626
rect 13014 13574 13020 13626
rect 13044 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13100 13626
rect 13124 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13180 13626
rect 13204 13574 13206 13626
rect 13206 13574 13258 13626
rect 13258 13574 13260 13626
rect 12884 13572 12940 13574
rect 12964 13572 13020 13574
rect 13044 13572 13100 13574
rect 13124 13572 13180 13574
rect 13204 13572 13260 13574
rect 7624 13082 7680 13084
rect 7704 13082 7760 13084
rect 7784 13082 7840 13084
rect 7864 13082 7920 13084
rect 7944 13082 8000 13084
rect 7624 13030 7626 13082
rect 7626 13030 7678 13082
rect 7678 13030 7680 13082
rect 7704 13030 7742 13082
rect 7742 13030 7754 13082
rect 7754 13030 7760 13082
rect 7784 13030 7806 13082
rect 7806 13030 7818 13082
rect 7818 13030 7840 13082
rect 7864 13030 7870 13082
rect 7870 13030 7882 13082
rect 7882 13030 7920 13082
rect 7944 13030 7946 13082
rect 7946 13030 7998 13082
rect 7998 13030 8000 13082
rect 7624 13028 7680 13030
rect 7704 13028 7760 13030
rect 7784 13028 7840 13030
rect 7864 13028 7920 13030
rect 7944 13028 8000 13030
rect 13624 13082 13680 13084
rect 13704 13082 13760 13084
rect 13784 13082 13840 13084
rect 13864 13082 13920 13084
rect 13944 13082 14000 13084
rect 13624 13030 13626 13082
rect 13626 13030 13678 13082
rect 13678 13030 13680 13082
rect 13704 13030 13742 13082
rect 13742 13030 13754 13082
rect 13754 13030 13760 13082
rect 13784 13030 13806 13082
rect 13806 13030 13818 13082
rect 13818 13030 13840 13082
rect 13864 13030 13870 13082
rect 13870 13030 13882 13082
rect 13882 13030 13920 13082
rect 13944 13030 13946 13082
rect 13946 13030 13998 13082
rect 13998 13030 14000 13082
rect 13624 13028 13680 13030
rect 13704 13028 13760 13030
rect 13784 13028 13840 13030
rect 13864 13028 13920 13030
rect 13944 13028 14000 13030
rect 6884 12538 6940 12540
rect 6964 12538 7020 12540
rect 7044 12538 7100 12540
rect 7124 12538 7180 12540
rect 7204 12538 7260 12540
rect 6884 12486 6886 12538
rect 6886 12486 6938 12538
rect 6938 12486 6940 12538
rect 6964 12486 7002 12538
rect 7002 12486 7014 12538
rect 7014 12486 7020 12538
rect 7044 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7100 12538
rect 7124 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7180 12538
rect 7204 12486 7206 12538
rect 7206 12486 7258 12538
rect 7258 12486 7260 12538
rect 6884 12484 6940 12486
rect 6964 12484 7020 12486
rect 7044 12484 7100 12486
rect 7124 12484 7180 12486
rect 7204 12484 7260 12486
rect 12884 12538 12940 12540
rect 12964 12538 13020 12540
rect 13044 12538 13100 12540
rect 13124 12538 13180 12540
rect 13204 12538 13260 12540
rect 12884 12486 12886 12538
rect 12886 12486 12938 12538
rect 12938 12486 12940 12538
rect 12964 12486 13002 12538
rect 13002 12486 13014 12538
rect 13014 12486 13020 12538
rect 13044 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13100 12538
rect 13124 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13180 12538
rect 13204 12486 13206 12538
rect 13206 12486 13258 12538
rect 13258 12486 13260 12538
rect 12884 12484 12940 12486
rect 12964 12484 13020 12486
rect 13044 12484 13100 12486
rect 13124 12484 13180 12486
rect 13204 12484 13260 12486
rect 7624 11994 7680 11996
rect 7704 11994 7760 11996
rect 7784 11994 7840 11996
rect 7864 11994 7920 11996
rect 7944 11994 8000 11996
rect 7624 11942 7626 11994
rect 7626 11942 7678 11994
rect 7678 11942 7680 11994
rect 7704 11942 7742 11994
rect 7742 11942 7754 11994
rect 7754 11942 7760 11994
rect 7784 11942 7806 11994
rect 7806 11942 7818 11994
rect 7818 11942 7840 11994
rect 7864 11942 7870 11994
rect 7870 11942 7882 11994
rect 7882 11942 7920 11994
rect 7944 11942 7946 11994
rect 7946 11942 7998 11994
rect 7998 11942 8000 11994
rect 7624 11940 7680 11942
rect 7704 11940 7760 11942
rect 7784 11940 7840 11942
rect 7864 11940 7920 11942
rect 7944 11940 8000 11942
rect 13624 11994 13680 11996
rect 13704 11994 13760 11996
rect 13784 11994 13840 11996
rect 13864 11994 13920 11996
rect 13944 11994 14000 11996
rect 13624 11942 13626 11994
rect 13626 11942 13678 11994
rect 13678 11942 13680 11994
rect 13704 11942 13742 11994
rect 13742 11942 13754 11994
rect 13754 11942 13760 11994
rect 13784 11942 13806 11994
rect 13806 11942 13818 11994
rect 13818 11942 13840 11994
rect 13864 11942 13870 11994
rect 13870 11942 13882 11994
rect 13882 11942 13920 11994
rect 13944 11942 13946 11994
rect 13946 11942 13998 11994
rect 13998 11942 14000 11994
rect 13624 11940 13680 11942
rect 13704 11940 13760 11942
rect 13784 11940 13840 11942
rect 13864 11940 13920 11942
rect 13944 11940 14000 11942
rect 6884 11450 6940 11452
rect 6964 11450 7020 11452
rect 7044 11450 7100 11452
rect 7124 11450 7180 11452
rect 7204 11450 7260 11452
rect 6884 11398 6886 11450
rect 6886 11398 6938 11450
rect 6938 11398 6940 11450
rect 6964 11398 7002 11450
rect 7002 11398 7014 11450
rect 7014 11398 7020 11450
rect 7044 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7100 11450
rect 7124 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7180 11450
rect 7204 11398 7206 11450
rect 7206 11398 7258 11450
rect 7258 11398 7260 11450
rect 6884 11396 6940 11398
rect 6964 11396 7020 11398
rect 7044 11396 7100 11398
rect 7124 11396 7180 11398
rect 7204 11396 7260 11398
rect 12884 11450 12940 11452
rect 12964 11450 13020 11452
rect 13044 11450 13100 11452
rect 13124 11450 13180 11452
rect 13204 11450 13260 11452
rect 12884 11398 12886 11450
rect 12886 11398 12938 11450
rect 12938 11398 12940 11450
rect 12964 11398 13002 11450
rect 13002 11398 13014 11450
rect 13014 11398 13020 11450
rect 13044 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13100 11450
rect 13124 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13180 11450
rect 13204 11398 13206 11450
rect 13206 11398 13258 11450
rect 13258 11398 13260 11450
rect 12884 11396 12940 11398
rect 12964 11396 13020 11398
rect 13044 11396 13100 11398
rect 13124 11396 13180 11398
rect 13204 11396 13260 11398
rect 7624 10906 7680 10908
rect 7704 10906 7760 10908
rect 7784 10906 7840 10908
rect 7864 10906 7920 10908
rect 7944 10906 8000 10908
rect 7624 10854 7626 10906
rect 7626 10854 7678 10906
rect 7678 10854 7680 10906
rect 7704 10854 7742 10906
rect 7742 10854 7754 10906
rect 7754 10854 7760 10906
rect 7784 10854 7806 10906
rect 7806 10854 7818 10906
rect 7818 10854 7840 10906
rect 7864 10854 7870 10906
rect 7870 10854 7882 10906
rect 7882 10854 7920 10906
rect 7944 10854 7946 10906
rect 7946 10854 7998 10906
rect 7998 10854 8000 10906
rect 7624 10852 7680 10854
rect 7704 10852 7760 10854
rect 7784 10852 7840 10854
rect 7864 10852 7920 10854
rect 7944 10852 8000 10854
rect 13624 10906 13680 10908
rect 13704 10906 13760 10908
rect 13784 10906 13840 10908
rect 13864 10906 13920 10908
rect 13944 10906 14000 10908
rect 13624 10854 13626 10906
rect 13626 10854 13678 10906
rect 13678 10854 13680 10906
rect 13704 10854 13742 10906
rect 13742 10854 13754 10906
rect 13754 10854 13760 10906
rect 13784 10854 13806 10906
rect 13806 10854 13818 10906
rect 13818 10854 13840 10906
rect 13864 10854 13870 10906
rect 13870 10854 13882 10906
rect 13882 10854 13920 10906
rect 13944 10854 13946 10906
rect 13946 10854 13998 10906
rect 13998 10854 14000 10906
rect 13624 10852 13680 10854
rect 13704 10852 13760 10854
rect 13784 10852 13840 10854
rect 13864 10852 13920 10854
rect 13944 10852 14000 10854
rect 6366 10240 6422 10296
rect 6884 10362 6940 10364
rect 6964 10362 7020 10364
rect 7044 10362 7100 10364
rect 7124 10362 7180 10364
rect 7204 10362 7260 10364
rect 6884 10310 6886 10362
rect 6886 10310 6938 10362
rect 6938 10310 6940 10362
rect 6964 10310 7002 10362
rect 7002 10310 7014 10362
rect 7014 10310 7020 10362
rect 7044 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7100 10362
rect 7124 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7180 10362
rect 7204 10310 7206 10362
rect 7206 10310 7258 10362
rect 7258 10310 7260 10362
rect 6884 10308 6940 10310
rect 6964 10308 7020 10310
rect 7044 10308 7100 10310
rect 7124 10308 7180 10310
rect 7204 10308 7260 10310
rect 12884 10362 12940 10364
rect 12964 10362 13020 10364
rect 13044 10362 13100 10364
rect 13124 10362 13180 10364
rect 13204 10362 13260 10364
rect 12884 10310 12886 10362
rect 12886 10310 12938 10362
rect 12938 10310 12940 10362
rect 12964 10310 13002 10362
rect 13002 10310 13014 10362
rect 13014 10310 13020 10362
rect 13044 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13100 10362
rect 13124 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13180 10362
rect 13204 10310 13206 10362
rect 13206 10310 13258 10362
rect 13258 10310 13260 10362
rect 12884 10308 12940 10310
rect 12964 10308 13020 10310
rect 13044 10308 13100 10310
rect 13124 10308 13180 10310
rect 13204 10308 13260 10310
rect 15198 10240 15254 10296
rect 4802 9560 4858 9616
rect 7624 9818 7680 9820
rect 7704 9818 7760 9820
rect 7784 9818 7840 9820
rect 7864 9818 7920 9820
rect 7944 9818 8000 9820
rect 7624 9766 7626 9818
rect 7626 9766 7678 9818
rect 7678 9766 7680 9818
rect 7704 9766 7742 9818
rect 7742 9766 7754 9818
rect 7754 9766 7760 9818
rect 7784 9766 7806 9818
rect 7806 9766 7818 9818
rect 7818 9766 7840 9818
rect 7864 9766 7870 9818
rect 7870 9766 7882 9818
rect 7882 9766 7920 9818
rect 7944 9766 7946 9818
rect 7946 9766 7998 9818
rect 7998 9766 8000 9818
rect 7624 9764 7680 9766
rect 7704 9764 7760 9766
rect 7784 9764 7840 9766
rect 7864 9764 7920 9766
rect 7944 9764 8000 9766
rect 13624 9818 13680 9820
rect 13704 9818 13760 9820
rect 13784 9818 13840 9820
rect 13864 9818 13920 9820
rect 13944 9818 14000 9820
rect 13624 9766 13626 9818
rect 13626 9766 13678 9818
rect 13678 9766 13680 9818
rect 13704 9766 13742 9818
rect 13742 9766 13754 9818
rect 13754 9766 13760 9818
rect 13784 9766 13806 9818
rect 13806 9766 13818 9818
rect 13818 9766 13840 9818
rect 13864 9766 13870 9818
rect 13870 9766 13882 9818
rect 13882 9766 13920 9818
rect 13944 9766 13946 9818
rect 13946 9766 13998 9818
rect 13998 9766 14000 9818
rect 13624 9764 13680 9766
rect 13704 9764 13760 9766
rect 13784 9764 13840 9766
rect 13864 9764 13920 9766
rect 13944 9764 14000 9766
rect 6884 9274 6940 9276
rect 6964 9274 7020 9276
rect 7044 9274 7100 9276
rect 7124 9274 7180 9276
rect 7204 9274 7260 9276
rect 6884 9222 6886 9274
rect 6886 9222 6938 9274
rect 6938 9222 6940 9274
rect 6964 9222 7002 9274
rect 7002 9222 7014 9274
rect 7014 9222 7020 9274
rect 7044 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7100 9274
rect 7124 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7180 9274
rect 7204 9222 7206 9274
rect 7206 9222 7258 9274
rect 7258 9222 7260 9274
rect 6884 9220 6940 9222
rect 6964 9220 7020 9222
rect 7044 9220 7100 9222
rect 7124 9220 7180 9222
rect 7204 9220 7260 9222
rect 12884 9274 12940 9276
rect 12964 9274 13020 9276
rect 13044 9274 13100 9276
rect 13124 9274 13180 9276
rect 13204 9274 13260 9276
rect 12884 9222 12886 9274
rect 12886 9222 12938 9274
rect 12938 9222 12940 9274
rect 12964 9222 13002 9274
rect 13002 9222 13014 9274
rect 13014 9222 13020 9274
rect 13044 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13100 9274
rect 13124 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13180 9274
rect 13204 9222 13206 9274
rect 13206 9222 13258 9274
rect 13258 9222 13260 9274
rect 12884 9220 12940 9222
rect 12964 9220 13020 9222
rect 13044 9220 13100 9222
rect 13124 9220 13180 9222
rect 13204 9220 13260 9222
rect 7624 8730 7680 8732
rect 7704 8730 7760 8732
rect 7784 8730 7840 8732
rect 7864 8730 7920 8732
rect 7944 8730 8000 8732
rect 7624 8678 7626 8730
rect 7626 8678 7678 8730
rect 7678 8678 7680 8730
rect 7704 8678 7742 8730
rect 7742 8678 7754 8730
rect 7754 8678 7760 8730
rect 7784 8678 7806 8730
rect 7806 8678 7818 8730
rect 7818 8678 7840 8730
rect 7864 8678 7870 8730
rect 7870 8678 7882 8730
rect 7882 8678 7920 8730
rect 7944 8678 7946 8730
rect 7946 8678 7998 8730
rect 7998 8678 8000 8730
rect 7624 8676 7680 8678
rect 7704 8676 7760 8678
rect 7784 8676 7840 8678
rect 7864 8676 7920 8678
rect 7944 8676 8000 8678
rect 13624 8730 13680 8732
rect 13704 8730 13760 8732
rect 13784 8730 13840 8732
rect 13864 8730 13920 8732
rect 13944 8730 14000 8732
rect 13624 8678 13626 8730
rect 13626 8678 13678 8730
rect 13678 8678 13680 8730
rect 13704 8678 13742 8730
rect 13742 8678 13754 8730
rect 13754 8678 13760 8730
rect 13784 8678 13806 8730
rect 13806 8678 13818 8730
rect 13818 8678 13840 8730
rect 13864 8678 13870 8730
rect 13870 8678 13882 8730
rect 13882 8678 13920 8730
rect 13944 8678 13946 8730
rect 13946 8678 13998 8730
rect 13998 8678 14000 8730
rect 13624 8676 13680 8678
rect 13704 8676 13760 8678
rect 13784 8676 13840 8678
rect 13864 8676 13920 8678
rect 13944 8676 14000 8678
rect 6884 8186 6940 8188
rect 6964 8186 7020 8188
rect 7044 8186 7100 8188
rect 7124 8186 7180 8188
rect 7204 8186 7260 8188
rect 6884 8134 6886 8186
rect 6886 8134 6938 8186
rect 6938 8134 6940 8186
rect 6964 8134 7002 8186
rect 7002 8134 7014 8186
rect 7014 8134 7020 8186
rect 7044 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7100 8186
rect 7124 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7180 8186
rect 7204 8134 7206 8186
rect 7206 8134 7258 8186
rect 7258 8134 7260 8186
rect 6884 8132 6940 8134
rect 6964 8132 7020 8134
rect 7044 8132 7100 8134
rect 7124 8132 7180 8134
rect 7204 8132 7260 8134
rect 12884 8186 12940 8188
rect 12964 8186 13020 8188
rect 13044 8186 13100 8188
rect 13124 8186 13180 8188
rect 13204 8186 13260 8188
rect 12884 8134 12886 8186
rect 12886 8134 12938 8186
rect 12938 8134 12940 8186
rect 12964 8134 13002 8186
rect 13002 8134 13014 8186
rect 13014 8134 13020 8186
rect 13044 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13100 8186
rect 13124 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13180 8186
rect 13204 8134 13206 8186
rect 13206 8134 13258 8186
rect 13258 8134 13260 8186
rect 12884 8132 12940 8134
rect 12964 8132 13020 8134
rect 13044 8132 13100 8134
rect 13124 8132 13180 8134
rect 13204 8132 13260 8134
rect 7624 7642 7680 7644
rect 7704 7642 7760 7644
rect 7784 7642 7840 7644
rect 7864 7642 7920 7644
rect 7944 7642 8000 7644
rect 7624 7590 7626 7642
rect 7626 7590 7678 7642
rect 7678 7590 7680 7642
rect 7704 7590 7742 7642
rect 7742 7590 7754 7642
rect 7754 7590 7760 7642
rect 7784 7590 7806 7642
rect 7806 7590 7818 7642
rect 7818 7590 7840 7642
rect 7864 7590 7870 7642
rect 7870 7590 7882 7642
rect 7882 7590 7920 7642
rect 7944 7590 7946 7642
rect 7946 7590 7998 7642
rect 7998 7590 8000 7642
rect 7624 7588 7680 7590
rect 7704 7588 7760 7590
rect 7784 7588 7840 7590
rect 7864 7588 7920 7590
rect 7944 7588 8000 7590
rect 13624 7642 13680 7644
rect 13704 7642 13760 7644
rect 13784 7642 13840 7644
rect 13864 7642 13920 7644
rect 13944 7642 14000 7644
rect 13624 7590 13626 7642
rect 13626 7590 13678 7642
rect 13678 7590 13680 7642
rect 13704 7590 13742 7642
rect 13742 7590 13754 7642
rect 13754 7590 13760 7642
rect 13784 7590 13806 7642
rect 13806 7590 13818 7642
rect 13818 7590 13840 7642
rect 13864 7590 13870 7642
rect 13870 7590 13882 7642
rect 13882 7590 13920 7642
rect 13944 7590 13946 7642
rect 13946 7590 13998 7642
rect 13998 7590 14000 7642
rect 13624 7588 13680 7590
rect 13704 7588 13760 7590
rect 13784 7588 13840 7590
rect 13864 7588 13920 7590
rect 13944 7588 14000 7590
rect 6884 7098 6940 7100
rect 6964 7098 7020 7100
rect 7044 7098 7100 7100
rect 7124 7098 7180 7100
rect 7204 7098 7260 7100
rect 6884 7046 6886 7098
rect 6886 7046 6938 7098
rect 6938 7046 6940 7098
rect 6964 7046 7002 7098
rect 7002 7046 7014 7098
rect 7014 7046 7020 7098
rect 7044 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7100 7098
rect 7124 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7180 7098
rect 7204 7046 7206 7098
rect 7206 7046 7258 7098
rect 7258 7046 7260 7098
rect 6884 7044 6940 7046
rect 6964 7044 7020 7046
rect 7044 7044 7100 7046
rect 7124 7044 7180 7046
rect 7204 7044 7260 7046
rect 12884 7098 12940 7100
rect 12964 7098 13020 7100
rect 13044 7098 13100 7100
rect 13124 7098 13180 7100
rect 13204 7098 13260 7100
rect 12884 7046 12886 7098
rect 12886 7046 12938 7098
rect 12938 7046 12940 7098
rect 12964 7046 13002 7098
rect 13002 7046 13014 7098
rect 13014 7046 13020 7098
rect 13044 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13100 7098
rect 13124 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13180 7098
rect 13204 7046 13206 7098
rect 13206 7046 13258 7098
rect 13258 7046 13260 7098
rect 12884 7044 12940 7046
rect 12964 7044 13020 7046
rect 13044 7044 13100 7046
rect 13124 7044 13180 7046
rect 13204 7044 13260 7046
rect 7624 6554 7680 6556
rect 7704 6554 7760 6556
rect 7784 6554 7840 6556
rect 7864 6554 7920 6556
rect 7944 6554 8000 6556
rect 7624 6502 7626 6554
rect 7626 6502 7678 6554
rect 7678 6502 7680 6554
rect 7704 6502 7742 6554
rect 7742 6502 7754 6554
rect 7754 6502 7760 6554
rect 7784 6502 7806 6554
rect 7806 6502 7818 6554
rect 7818 6502 7840 6554
rect 7864 6502 7870 6554
rect 7870 6502 7882 6554
rect 7882 6502 7920 6554
rect 7944 6502 7946 6554
rect 7946 6502 7998 6554
rect 7998 6502 8000 6554
rect 7624 6500 7680 6502
rect 7704 6500 7760 6502
rect 7784 6500 7840 6502
rect 7864 6500 7920 6502
rect 7944 6500 8000 6502
rect 13624 6554 13680 6556
rect 13704 6554 13760 6556
rect 13784 6554 13840 6556
rect 13864 6554 13920 6556
rect 13944 6554 14000 6556
rect 13624 6502 13626 6554
rect 13626 6502 13678 6554
rect 13678 6502 13680 6554
rect 13704 6502 13742 6554
rect 13742 6502 13754 6554
rect 13754 6502 13760 6554
rect 13784 6502 13806 6554
rect 13806 6502 13818 6554
rect 13818 6502 13840 6554
rect 13864 6502 13870 6554
rect 13870 6502 13882 6554
rect 13882 6502 13920 6554
rect 13944 6502 13946 6554
rect 13946 6502 13998 6554
rect 13998 6502 14000 6554
rect 13624 6500 13680 6502
rect 13704 6500 13760 6502
rect 13784 6500 13840 6502
rect 13864 6500 13920 6502
rect 13944 6500 14000 6502
<< metal3 >>
rect 6874 13632 7270 13633
rect 6874 13568 6880 13632
rect 6944 13568 6960 13632
rect 7024 13568 7040 13632
rect 7104 13568 7120 13632
rect 7184 13568 7200 13632
rect 7264 13568 7270 13632
rect 6874 13567 7270 13568
rect 12874 13632 13270 13633
rect 12874 13568 12880 13632
rect 12944 13568 12960 13632
rect 13024 13568 13040 13632
rect 13104 13568 13120 13632
rect 13184 13568 13200 13632
rect 13264 13568 13270 13632
rect 12874 13567 13270 13568
rect 7614 13088 8010 13089
rect 7614 13024 7620 13088
rect 7684 13024 7700 13088
rect 7764 13024 7780 13088
rect 7844 13024 7860 13088
rect 7924 13024 7940 13088
rect 8004 13024 8010 13088
rect 7614 13023 8010 13024
rect 13614 13088 14010 13089
rect 13614 13024 13620 13088
rect 13684 13024 13700 13088
rect 13764 13024 13780 13088
rect 13844 13024 13860 13088
rect 13924 13024 13940 13088
rect 14004 13024 14010 13088
rect 13614 13023 14010 13024
rect 6874 12544 7270 12545
rect 6874 12480 6880 12544
rect 6944 12480 6960 12544
rect 7024 12480 7040 12544
rect 7104 12480 7120 12544
rect 7184 12480 7200 12544
rect 7264 12480 7270 12544
rect 6874 12479 7270 12480
rect 12874 12544 13270 12545
rect 12874 12480 12880 12544
rect 12944 12480 12960 12544
rect 13024 12480 13040 12544
rect 13104 12480 13120 12544
rect 13184 12480 13200 12544
rect 13264 12480 13270 12544
rect 12874 12479 13270 12480
rect 7614 12000 8010 12001
rect 7614 11936 7620 12000
rect 7684 11936 7700 12000
rect 7764 11936 7780 12000
rect 7844 11936 7860 12000
rect 7924 11936 7940 12000
rect 8004 11936 8010 12000
rect 7614 11935 8010 11936
rect 13614 12000 14010 12001
rect 13614 11936 13620 12000
rect 13684 11936 13700 12000
rect 13764 11936 13780 12000
rect 13844 11936 13860 12000
rect 13924 11936 13940 12000
rect 14004 11936 14010 12000
rect 13614 11935 14010 11936
rect 6874 11456 7270 11457
rect 6874 11392 6880 11456
rect 6944 11392 6960 11456
rect 7024 11392 7040 11456
rect 7104 11392 7120 11456
rect 7184 11392 7200 11456
rect 7264 11392 7270 11456
rect 6874 11391 7270 11392
rect 12874 11456 13270 11457
rect 12874 11392 12880 11456
rect 12944 11392 12960 11456
rect 13024 11392 13040 11456
rect 13104 11392 13120 11456
rect 13184 11392 13200 11456
rect 13264 11392 13270 11456
rect 12874 11391 13270 11392
rect 7614 10912 8010 10913
rect 7614 10848 7620 10912
rect 7684 10848 7700 10912
rect 7764 10848 7780 10912
rect 7844 10848 7860 10912
rect 7924 10848 7940 10912
rect 8004 10848 8010 10912
rect 7614 10847 8010 10848
rect 13614 10912 14010 10913
rect 13614 10848 13620 10912
rect 13684 10848 13700 10912
rect 13764 10848 13780 10912
rect 13844 10848 13860 10912
rect 13924 10848 13940 10912
rect 14004 10848 14010 10912
rect 13614 10847 14010 10848
rect 6874 10368 7270 10369
rect 0 10298 800 10328
rect 6874 10304 6880 10368
rect 6944 10304 6960 10368
rect 7024 10304 7040 10368
rect 7104 10304 7120 10368
rect 7184 10304 7200 10368
rect 7264 10304 7270 10368
rect 6874 10303 7270 10304
rect 12874 10368 13270 10369
rect 12874 10304 12880 10368
rect 12944 10304 12960 10368
rect 13024 10304 13040 10368
rect 13104 10304 13120 10368
rect 13184 10304 13200 10368
rect 13264 10304 13270 10368
rect 12874 10303 13270 10304
rect 6361 10298 6427 10301
rect 0 10296 6427 10298
rect 0 10240 6366 10296
rect 6422 10240 6427 10296
rect 0 10238 6427 10240
rect 0 10208 800 10238
rect 6361 10235 6427 10238
rect 15193 10298 15259 10301
rect 19200 10298 20000 10328
rect 15193 10296 20000 10298
rect 15193 10240 15198 10296
rect 15254 10240 20000 10296
rect 15193 10238 20000 10240
rect 15193 10235 15259 10238
rect 19200 10208 20000 10238
rect 7614 9824 8010 9825
rect 7614 9760 7620 9824
rect 7684 9760 7700 9824
rect 7764 9760 7780 9824
rect 7844 9760 7860 9824
rect 7924 9760 7940 9824
rect 8004 9760 8010 9824
rect 7614 9759 8010 9760
rect 13614 9824 14010 9825
rect 13614 9760 13620 9824
rect 13684 9760 13700 9824
rect 13764 9760 13780 9824
rect 13844 9760 13860 9824
rect 13924 9760 13940 9824
rect 14004 9760 14010 9824
rect 13614 9759 14010 9760
rect 0 9618 800 9648
rect 4797 9618 4863 9621
rect 0 9616 4863 9618
rect 0 9560 4802 9616
rect 4858 9560 4863 9616
rect 0 9558 4863 9560
rect 0 9528 800 9558
rect 4797 9555 4863 9558
rect 6874 9280 7270 9281
rect 6874 9216 6880 9280
rect 6944 9216 6960 9280
rect 7024 9216 7040 9280
rect 7104 9216 7120 9280
rect 7184 9216 7200 9280
rect 7264 9216 7270 9280
rect 6874 9215 7270 9216
rect 12874 9280 13270 9281
rect 12874 9216 12880 9280
rect 12944 9216 12960 9280
rect 13024 9216 13040 9280
rect 13104 9216 13120 9280
rect 13184 9216 13200 9280
rect 13264 9216 13270 9280
rect 12874 9215 13270 9216
rect 7614 8736 8010 8737
rect 7614 8672 7620 8736
rect 7684 8672 7700 8736
rect 7764 8672 7780 8736
rect 7844 8672 7860 8736
rect 7924 8672 7940 8736
rect 8004 8672 8010 8736
rect 7614 8671 8010 8672
rect 13614 8736 14010 8737
rect 13614 8672 13620 8736
rect 13684 8672 13700 8736
rect 13764 8672 13780 8736
rect 13844 8672 13860 8736
rect 13924 8672 13940 8736
rect 14004 8672 14010 8736
rect 13614 8671 14010 8672
rect 6874 8192 7270 8193
rect 6874 8128 6880 8192
rect 6944 8128 6960 8192
rect 7024 8128 7040 8192
rect 7104 8128 7120 8192
rect 7184 8128 7200 8192
rect 7264 8128 7270 8192
rect 6874 8127 7270 8128
rect 12874 8192 13270 8193
rect 12874 8128 12880 8192
rect 12944 8128 12960 8192
rect 13024 8128 13040 8192
rect 13104 8128 13120 8192
rect 13184 8128 13200 8192
rect 13264 8128 13270 8192
rect 12874 8127 13270 8128
rect 7614 7648 8010 7649
rect 7614 7584 7620 7648
rect 7684 7584 7700 7648
rect 7764 7584 7780 7648
rect 7844 7584 7860 7648
rect 7924 7584 7940 7648
rect 8004 7584 8010 7648
rect 7614 7583 8010 7584
rect 13614 7648 14010 7649
rect 13614 7584 13620 7648
rect 13684 7584 13700 7648
rect 13764 7584 13780 7648
rect 13844 7584 13860 7648
rect 13924 7584 13940 7648
rect 14004 7584 14010 7648
rect 13614 7583 14010 7584
rect 6874 7104 7270 7105
rect 6874 7040 6880 7104
rect 6944 7040 6960 7104
rect 7024 7040 7040 7104
rect 7104 7040 7120 7104
rect 7184 7040 7200 7104
rect 7264 7040 7270 7104
rect 6874 7039 7270 7040
rect 12874 7104 13270 7105
rect 12874 7040 12880 7104
rect 12944 7040 12960 7104
rect 13024 7040 13040 7104
rect 13104 7040 13120 7104
rect 13184 7040 13200 7104
rect 13264 7040 13270 7104
rect 12874 7039 13270 7040
rect 7614 6560 8010 6561
rect 7614 6496 7620 6560
rect 7684 6496 7700 6560
rect 7764 6496 7780 6560
rect 7844 6496 7860 6560
rect 7924 6496 7940 6560
rect 8004 6496 8010 6560
rect 7614 6495 8010 6496
rect 13614 6560 14010 6561
rect 13614 6496 13620 6560
rect 13684 6496 13700 6560
rect 13764 6496 13780 6560
rect 13844 6496 13860 6560
rect 13924 6496 13940 6560
rect 14004 6496 14010 6560
rect 13614 6495 14010 6496
<< via3 >>
rect 6880 13628 6944 13632
rect 6880 13572 6884 13628
rect 6884 13572 6940 13628
rect 6940 13572 6944 13628
rect 6880 13568 6944 13572
rect 6960 13628 7024 13632
rect 6960 13572 6964 13628
rect 6964 13572 7020 13628
rect 7020 13572 7024 13628
rect 6960 13568 7024 13572
rect 7040 13628 7104 13632
rect 7040 13572 7044 13628
rect 7044 13572 7100 13628
rect 7100 13572 7104 13628
rect 7040 13568 7104 13572
rect 7120 13628 7184 13632
rect 7120 13572 7124 13628
rect 7124 13572 7180 13628
rect 7180 13572 7184 13628
rect 7120 13568 7184 13572
rect 7200 13628 7264 13632
rect 7200 13572 7204 13628
rect 7204 13572 7260 13628
rect 7260 13572 7264 13628
rect 7200 13568 7264 13572
rect 12880 13628 12944 13632
rect 12880 13572 12884 13628
rect 12884 13572 12940 13628
rect 12940 13572 12944 13628
rect 12880 13568 12944 13572
rect 12960 13628 13024 13632
rect 12960 13572 12964 13628
rect 12964 13572 13020 13628
rect 13020 13572 13024 13628
rect 12960 13568 13024 13572
rect 13040 13628 13104 13632
rect 13040 13572 13044 13628
rect 13044 13572 13100 13628
rect 13100 13572 13104 13628
rect 13040 13568 13104 13572
rect 13120 13628 13184 13632
rect 13120 13572 13124 13628
rect 13124 13572 13180 13628
rect 13180 13572 13184 13628
rect 13120 13568 13184 13572
rect 13200 13628 13264 13632
rect 13200 13572 13204 13628
rect 13204 13572 13260 13628
rect 13260 13572 13264 13628
rect 13200 13568 13264 13572
rect 7620 13084 7684 13088
rect 7620 13028 7624 13084
rect 7624 13028 7680 13084
rect 7680 13028 7684 13084
rect 7620 13024 7684 13028
rect 7700 13084 7764 13088
rect 7700 13028 7704 13084
rect 7704 13028 7760 13084
rect 7760 13028 7764 13084
rect 7700 13024 7764 13028
rect 7780 13084 7844 13088
rect 7780 13028 7784 13084
rect 7784 13028 7840 13084
rect 7840 13028 7844 13084
rect 7780 13024 7844 13028
rect 7860 13084 7924 13088
rect 7860 13028 7864 13084
rect 7864 13028 7920 13084
rect 7920 13028 7924 13084
rect 7860 13024 7924 13028
rect 7940 13084 8004 13088
rect 7940 13028 7944 13084
rect 7944 13028 8000 13084
rect 8000 13028 8004 13084
rect 7940 13024 8004 13028
rect 13620 13084 13684 13088
rect 13620 13028 13624 13084
rect 13624 13028 13680 13084
rect 13680 13028 13684 13084
rect 13620 13024 13684 13028
rect 13700 13084 13764 13088
rect 13700 13028 13704 13084
rect 13704 13028 13760 13084
rect 13760 13028 13764 13084
rect 13700 13024 13764 13028
rect 13780 13084 13844 13088
rect 13780 13028 13784 13084
rect 13784 13028 13840 13084
rect 13840 13028 13844 13084
rect 13780 13024 13844 13028
rect 13860 13084 13924 13088
rect 13860 13028 13864 13084
rect 13864 13028 13920 13084
rect 13920 13028 13924 13084
rect 13860 13024 13924 13028
rect 13940 13084 14004 13088
rect 13940 13028 13944 13084
rect 13944 13028 14000 13084
rect 14000 13028 14004 13084
rect 13940 13024 14004 13028
rect 6880 12540 6944 12544
rect 6880 12484 6884 12540
rect 6884 12484 6940 12540
rect 6940 12484 6944 12540
rect 6880 12480 6944 12484
rect 6960 12540 7024 12544
rect 6960 12484 6964 12540
rect 6964 12484 7020 12540
rect 7020 12484 7024 12540
rect 6960 12480 7024 12484
rect 7040 12540 7104 12544
rect 7040 12484 7044 12540
rect 7044 12484 7100 12540
rect 7100 12484 7104 12540
rect 7040 12480 7104 12484
rect 7120 12540 7184 12544
rect 7120 12484 7124 12540
rect 7124 12484 7180 12540
rect 7180 12484 7184 12540
rect 7120 12480 7184 12484
rect 7200 12540 7264 12544
rect 7200 12484 7204 12540
rect 7204 12484 7260 12540
rect 7260 12484 7264 12540
rect 7200 12480 7264 12484
rect 12880 12540 12944 12544
rect 12880 12484 12884 12540
rect 12884 12484 12940 12540
rect 12940 12484 12944 12540
rect 12880 12480 12944 12484
rect 12960 12540 13024 12544
rect 12960 12484 12964 12540
rect 12964 12484 13020 12540
rect 13020 12484 13024 12540
rect 12960 12480 13024 12484
rect 13040 12540 13104 12544
rect 13040 12484 13044 12540
rect 13044 12484 13100 12540
rect 13100 12484 13104 12540
rect 13040 12480 13104 12484
rect 13120 12540 13184 12544
rect 13120 12484 13124 12540
rect 13124 12484 13180 12540
rect 13180 12484 13184 12540
rect 13120 12480 13184 12484
rect 13200 12540 13264 12544
rect 13200 12484 13204 12540
rect 13204 12484 13260 12540
rect 13260 12484 13264 12540
rect 13200 12480 13264 12484
rect 7620 11996 7684 12000
rect 7620 11940 7624 11996
rect 7624 11940 7680 11996
rect 7680 11940 7684 11996
rect 7620 11936 7684 11940
rect 7700 11996 7764 12000
rect 7700 11940 7704 11996
rect 7704 11940 7760 11996
rect 7760 11940 7764 11996
rect 7700 11936 7764 11940
rect 7780 11996 7844 12000
rect 7780 11940 7784 11996
rect 7784 11940 7840 11996
rect 7840 11940 7844 11996
rect 7780 11936 7844 11940
rect 7860 11996 7924 12000
rect 7860 11940 7864 11996
rect 7864 11940 7920 11996
rect 7920 11940 7924 11996
rect 7860 11936 7924 11940
rect 7940 11996 8004 12000
rect 7940 11940 7944 11996
rect 7944 11940 8000 11996
rect 8000 11940 8004 11996
rect 7940 11936 8004 11940
rect 13620 11996 13684 12000
rect 13620 11940 13624 11996
rect 13624 11940 13680 11996
rect 13680 11940 13684 11996
rect 13620 11936 13684 11940
rect 13700 11996 13764 12000
rect 13700 11940 13704 11996
rect 13704 11940 13760 11996
rect 13760 11940 13764 11996
rect 13700 11936 13764 11940
rect 13780 11996 13844 12000
rect 13780 11940 13784 11996
rect 13784 11940 13840 11996
rect 13840 11940 13844 11996
rect 13780 11936 13844 11940
rect 13860 11996 13924 12000
rect 13860 11940 13864 11996
rect 13864 11940 13920 11996
rect 13920 11940 13924 11996
rect 13860 11936 13924 11940
rect 13940 11996 14004 12000
rect 13940 11940 13944 11996
rect 13944 11940 14000 11996
rect 14000 11940 14004 11996
rect 13940 11936 14004 11940
rect 6880 11452 6944 11456
rect 6880 11396 6884 11452
rect 6884 11396 6940 11452
rect 6940 11396 6944 11452
rect 6880 11392 6944 11396
rect 6960 11452 7024 11456
rect 6960 11396 6964 11452
rect 6964 11396 7020 11452
rect 7020 11396 7024 11452
rect 6960 11392 7024 11396
rect 7040 11452 7104 11456
rect 7040 11396 7044 11452
rect 7044 11396 7100 11452
rect 7100 11396 7104 11452
rect 7040 11392 7104 11396
rect 7120 11452 7184 11456
rect 7120 11396 7124 11452
rect 7124 11396 7180 11452
rect 7180 11396 7184 11452
rect 7120 11392 7184 11396
rect 7200 11452 7264 11456
rect 7200 11396 7204 11452
rect 7204 11396 7260 11452
rect 7260 11396 7264 11452
rect 7200 11392 7264 11396
rect 12880 11452 12944 11456
rect 12880 11396 12884 11452
rect 12884 11396 12940 11452
rect 12940 11396 12944 11452
rect 12880 11392 12944 11396
rect 12960 11452 13024 11456
rect 12960 11396 12964 11452
rect 12964 11396 13020 11452
rect 13020 11396 13024 11452
rect 12960 11392 13024 11396
rect 13040 11452 13104 11456
rect 13040 11396 13044 11452
rect 13044 11396 13100 11452
rect 13100 11396 13104 11452
rect 13040 11392 13104 11396
rect 13120 11452 13184 11456
rect 13120 11396 13124 11452
rect 13124 11396 13180 11452
rect 13180 11396 13184 11452
rect 13120 11392 13184 11396
rect 13200 11452 13264 11456
rect 13200 11396 13204 11452
rect 13204 11396 13260 11452
rect 13260 11396 13264 11452
rect 13200 11392 13264 11396
rect 7620 10908 7684 10912
rect 7620 10852 7624 10908
rect 7624 10852 7680 10908
rect 7680 10852 7684 10908
rect 7620 10848 7684 10852
rect 7700 10908 7764 10912
rect 7700 10852 7704 10908
rect 7704 10852 7760 10908
rect 7760 10852 7764 10908
rect 7700 10848 7764 10852
rect 7780 10908 7844 10912
rect 7780 10852 7784 10908
rect 7784 10852 7840 10908
rect 7840 10852 7844 10908
rect 7780 10848 7844 10852
rect 7860 10908 7924 10912
rect 7860 10852 7864 10908
rect 7864 10852 7920 10908
rect 7920 10852 7924 10908
rect 7860 10848 7924 10852
rect 7940 10908 8004 10912
rect 7940 10852 7944 10908
rect 7944 10852 8000 10908
rect 8000 10852 8004 10908
rect 7940 10848 8004 10852
rect 13620 10908 13684 10912
rect 13620 10852 13624 10908
rect 13624 10852 13680 10908
rect 13680 10852 13684 10908
rect 13620 10848 13684 10852
rect 13700 10908 13764 10912
rect 13700 10852 13704 10908
rect 13704 10852 13760 10908
rect 13760 10852 13764 10908
rect 13700 10848 13764 10852
rect 13780 10908 13844 10912
rect 13780 10852 13784 10908
rect 13784 10852 13840 10908
rect 13840 10852 13844 10908
rect 13780 10848 13844 10852
rect 13860 10908 13924 10912
rect 13860 10852 13864 10908
rect 13864 10852 13920 10908
rect 13920 10852 13924 10908
rect 13860 10848 13924 10852
rect 13940 10908 14004 10912
rect 13940 10852 13944 10908
rect 13944 10852 14000 10908
rect 14000 10852 14004 10908
rect 13940 10848 14004 10852
rect 6880 10364 6944 10368
rect 6880 10308 6884 10364
rect 6884 10308 6940 10364
rect 6940 10308 6944 10364
rect 6880 10304 6944 10308
rect 6960 10364 7024 10368
rect 6960 10308 6964 10364
rect 6964 10308 7020 10364
rect 7020 10308 7024 10364
rect 6960 10304 7024 10308
rect 7040 10364 7104 10368
rect 7040 10308 7044 10364
rect 7044 10308 7100 10364
rect 7100 10308 7104 10364
rect 7040 10304 7104 10308
rect 7120 10364 7184 10368
rect 7120 10308 7124 10364
rect 7124 10308 7180 10364
rect 7180 10308 7184 10364
rect 7120 10304 7184 10308
rect 7200 10364 7264 10368
rect 7200 10308 7204 10364
rect 7204 10308 7260 10364
rect 7260 10308 7264 10364
rect 7200 10304 7264 10308
rect 12880 10364 12944 10368
rect 12880 10308 12884 10364
rect 12884 10308 12940 10364
rect 12940 10308 12944 10364
rect 12880 10304 12944 10308
rect 12960 10364 13024 10368
rect 12960 10308 12964 10364
rect 12964 10308 13020 10364
rect 13020 10308 13024 10364
rect 12960 10304 13024 10308
rect 13040 10364 13104 10368
rect 13040 10308 13044 10364
rect 13044 10308 13100 10364
rect 13100 10308 13104 10364
rect 13040 10304 13104 10308
rect 13120 10364 13184 10368
rect 13120 10308 13124 10364
rect 13124 10308 13180 10364
rect 13180 10308 13184 10364
rect 13120 10304 13184 10308
rect 13200 10364 13264 10368
rect 13200 10308 13204 10364
rect 13204 10308 13260 10364
rect 13260 10308 13264 10364
rect 13200 10304 13264 10308
rect 7620 9820 7684 9824
rect 7620 9764 7624 9820
rect 7624 9764 7680 9820
rect 7680 9764 7684 9820
rect 7620 9760 7684 9764
rect 7700 9820 7764 9824
rect 7700 9764 7704 9820
rect 7704 9764 7760 9820
rect 7760 9764 7764 9820
rect 7700 9760 7764 9764
rect 7780 9820 7844 9824
rect 7780 9764 7784 9820
rect 7784 9764 7840 9820
rect 7840 9764 7844 9820
rect 7780 9760 7844 9764
rect 7860 9820 7924 9824
rect 7860 9764 7864 9820
rect 7864 9764 7920 9820
rect 7920 9764 7924 9820
rect 7860 9760 7924 9764
rect 7940 9820 8004 9824
rect 7940 9764 7944 9820
rect 7944 9764 8000 9820
rect 8000 9764 8004 9820
rect 7940 9760 8004 9764
rect 13620 9820 13684 9824
rect 13620 9764 13624 9820
rect 13624 9764 13680 9820
rect 13680 9764 13684 9820
rect 13620 9760 13684 9764
rect 13700 9820 13764 9824
rect 13700 9764 13704 9820
rect 13704 9764 13760 9820
rect 13760 9764 13764 9820
rect 13700 9760 13764 9764
rect 13780 9820 13844 9824
rect 13780 9764 13784 9820
rect 13784 9764 13840 9820
rect 13840 9764 13844 9820
rect 13780 9760 13844 9764
rect 13860 9820 13924 9824
rect 13860 9764 13864 9820
rect 13864 9764 13920 9820
rect 13920 9764 13924 9820
rect 13860 9760 13924 9764
rect 13940 9820 14004 9824
rect 13940 9764 13944 9820
rect 13944 9764 14000 9820
rect 14000 9764 14004 9820
rect 13940 9760 14004 9764
rect 6880 9276 6944 9280
rect 6880 9220 6884 9276
rect 6884 9220 6940 9276
rect 6940 9220 6944 9276
rect 6880 9216 6944 9220
rect 6960 9276 7024 9280
rect 6960 9220 6964 9276
rect 6964 9220 7020 9276
rect 7020 9220 7024 9276
rect 6960 9216 7024 9220
rect 7040 9276 7104 9280
rect 7040 9220 7044 9276
rect 7044 9220 7100 9276
rect 7100 9220 7104 9276
rect 7040 9216 7104 9220
rect 7120 9276 7184 9280
rect 7120 9220 7124 9276
rect 7124 9220 7180 9276
rect 7180 9220 7184 9276
rect 7120 9216 7184 9220
rect 7200 9276 7264 9280
rect 7200 9220 7204 9276
rect 7204 9220 7260 9276
rect 7260 9220 7264 9276
rect 7200 9216 7264 9220
rect 12880 9276 12944 9280
rect 12880 9220 12884 9276
rect 12884 9220 12940 9276
rect 12940 9220 12944 9276
rect 12880 9216 12944 9220
rect 12960 9276 13024 9280
rect 12960 9220 12964 9276
rect 12964 9220 13020 9276
rect 13020 9220 13024 9276
rect 12960 9216 13024 9220
rect 13040 9276 13104 9280
rect 13040 9220 13044 9276
rect 13044 9220 13100 9276
rect 13100 9220 13104 9276
rect 13040 9216 13104 9220
rect 13120 9276 13184 9280
rect 13120 9220 13124 9276
rect 13124 9220 13180 9276
rect 13180 9220 13184 9276
rect 13120 9216 13184 9220
rect 13200 9276 13264 9280
rect 13200 9220 13204 9276
rect 13204 9220 13260 9276
rect 13260 9220 13264 9276
rect 13200 9216 13264 9220
rect 7620 8732 7684 8736
rect 7620 8676 7624 8732
rect 7624 8676 7680 8732
rect 7680 8676 7684 8732
rect 7620 8672 7684 8676
rect 7700 8732 7764 8736
rect 7700 8676 7704 8732
rect 7704 8676 7760 8732
rect 7760 8676 7764 8732
rect 7700 8672 7764 8676
rect 7780 8732 7844 8736
rect 7780 8676 7784 8732
rect 7784 8676 7840 8732
rect 7840 8676 7844 8732
rect 7780 8672 7844 8676
rect 7860 8732 7924 8736
rect 7860 8676 7864 8732
rect 7864 8676 7920 8732
rect 7920 8676 7924 8732
rect 7860 8672 7924 8676
rect 7940 8732 8004 8736
rect 7940 8676 7944 8732
rect 7944 8676 8000 8732
rect 8000 8676 8004 8732
rect 7940 8672 8004 8676
rect 13620 8732 13684 8736
rect 13620 8676 13624 8732
rect 13624 8676 13680 8732
rect 13680 8676 13684 8732
rect 13620 8672 13684 8676
rect 13700 8732 13764 8736
rect 13700 8676 13704 8732
rect 13704 8676 13760 8732
rect 13760 8676 13764 8732
rect 13700 8672 13764 8676
rect 13780 8732 13844 8736
rect 13780 8676 13784 8732
rect 13784 8676 13840 8732
rect 13840 8676 13844 8732
rect 13780 8672 13844 8676
rect 13860 8732 13924 8736
rect 13860 8676 13864 8732
rect 13864 8676 13920 8732
rect 13920 8676 13924 8732
rect 13860 8672 13924 8676
rect 13940 8732 14004 8736
rect 13940 8676 13944 8732
rect 13944 8676 14000 8732
rect 14000 8676 14004 8732
rect 13940 8672 14004 8676
rect 6880 8188 6944 8192
rect 6880 8132 6884 8188
rect 6884 8132 6940 8188
rect 6940 8132 6944 8188
rect 6880 8128 6944 8132
rect 6960 8188 7024 8192
rect 6960 8132 6964 8188
rect 6964 8132 7020 8188
rect 7020 8132 7024 8188
rect 6960 8128 7024 8132
rect 7040 8188 7104 8192
rect 7040 8132 7044 8188
rect 7044 8132 7100 8188
rect 7100 8132 7104 8188
rect 7040 8128 7104 8132
rect 7120 8188 7184 8192
rect 7120 8132 7124 8188
rect 7124 8132 7180 8188
rect 7180 8132 7184 8188
rect 7120 8128 7184 8132
rect 7200 8188 7264 8192
rect 7200 8132 7204 8188
rect 7204 8132 7260 8188
rect 7260 8132 7264 8188
rect 7200 8128 7264 8132
rect 12880 8188 12944 8192
rect 12880 8132 12884 8188
rect 12884 8132 12940 8188
rect 12940 8132 12944 8188
rect 12880 8128 12944 8132
rect 12960 8188 13024 8192
rect 12960 8132 12964 8188
rect 12964 8132 13020 8188
rect 13020 8132 13024 8188
rect 12960 8128 13024 8132
rect 13040 8188 13104 8192
rect 13040 8132 13044 8188
rect 13044 8132 13100 8188
rect 13100 8132 13104 8188
rect 13040 8128 13104 8132
rect 13120 8188 13184 8192
rect 13120 8132 13124 8188
rect 13124 8132 13180 8188
rect 13180 8132 13184 8188
rect 13120 8128 13184 8132
rect 13200 8188 13264 8192
rect 13200 8132 13204 8188
rect 13204 8132 13260 8188
rect 13260 8132 13264 8188
rect 13200 8128 13264 8132
rect 7620 7644 7684 7648
rect 7620 7588 7624 7644
rect 7624 7588 7680 7644
rect 7680 7588 7684 7644
rect 7620 7584 7684 7588
rect 7700 7644 7764 7648
rect 7700 7588 7704 7644
rect 7704 7588 7760 7644
rect 7760 7588 7764 7644
rect 7700 7584 7764 7588
rect 7780 7644 7844 7648
rect 7780 7588 7784 7644
rect 7784 7588 7840 7644
rect 7840 7588 7844 7644
rect 7780 7584 7844 7588
rect 7860 7644 7924 7648
rect 7860 7588 7864 7644
rect 7864 7588 7920 7644
rect 7920 7588 7924 7644
rect 7860 7584 7924 7588
rect 7940 7644 8004 7648
rect 7940 7588 7944 7644
rect 7944 7588 8000 7644
rect 8000 7588 8004 7644
rect 7940 7584 8004 7588
rect 13620 7644 13684 7648
rect 13620 7588 13624 7644
rect 13624 7588 13680 7644
rect 13680 7588 13684 7644
rect 13620 7584 13684 7588
rect 13700 7644 13764 7648
rect 13700 7588 13704 7644
rect 13704 7588 13760 7644
rect 13760 7588 13764 7644
rect 13700 7584 13764 7588
rect 13780 7644 13844 7648
rect 13780 7588 13784 7644
rect 13784 7588 13840 7644
rect 13840 7588 13844 7644
rect 13780 7584 13844 7588
rect 13860 7644 13924 7648
rect 13860 7588 13864 7644
rect 13864 7588 13920 7644
rect 13920 7588 13924 7644
rect 13860 7584 13924 7588
rect 13940 7644 14004 7648
rect 13940 7588 13944 7644
rect 13944 7588 14000 7644
rect 14000 7588 14004 7644
rect 13940 7584 14004 7588
rect 6880 7100 6944 7104
rect 6880 7044 6884 7100
rect 6884 7044 6940 7100
rect 6940 7044 6944 7100
rect 6880 7040 6944 7044
rect 6960 7100 7024 7104
rect 6960 7044 6964 7100
rect 6964 7044 7020 7100
rect 7020 7044 7024 7100
rect 6960 7040 7024 7044
rect 7040 7100 7104 7104
rect 7040 7044 7044 7100
rect 7044 7044 7100 7100
rect 7100 7044 7104 7100
rect 7040 7040 7104 7044
rect 7120 7100 7184 7104
rect 7120 7044 7124 7100
rect 7124 7044 7180 7100
rect 7180 7044 7184 7100
rect 7120 7040 7184 7044
rect 7200 7100 7264 7104
rect 7200 7044 7204 7100
rect 7204 7044 7260 7100
rect 7260 7044 7264 7100
rect 7200 7040 7264 7044
rect 12880 7100 12944 7104
rect 12880 7044 12884 7100
rect 12884 7044 12940 7100
rect 12940 7044 12944 7100
rect 12880 7040 12944 7044
rect 12960 7100 13024 7104
rect 12960 7044 12964 7100
rect 12964 7044 13020 7100
rect 13020 7044 13024 7100
rect 12960 7040 13024 7044
rect 13040 7100 13104 7104
rect 13040 7044 13044 7100
rect 13044 7044 13100 7100
rect 13100 7044 13104 7100
rect 13040 7040 13104 7044
rect 13120 7100 13184 7104
rect 13120 7044 13124 7100
rect 13124 7044 13180 7100
rect 13180 7044 13184 7100
rect 13120 7040 13184 7044
rect 13200 7100 13264 7104
rect 13200 7044 13204 7100
rect 13204 7044 13260 7100
rect 13260 7044 13264 7100
rect 13200 7040 13264 7044
rect 7620 6556 7684 6560
rect 7620 6500 7624 6556
rect 7624 6500 7680 6556
rect 7680 6500 7684 6556
rect 7620 6496 7684 6500
rect 7700 6556 7764 6560
rect 7700 6500 7704 6556
rect 7704 6500 7760 6556
rect 7760 6500 7764 6556
rect 7700 6496 7764 6500
rect 7780 6556 7844 6560
rect 7780 6500 7784 6556
rect 7784 6500 7840 6556
rect 7840 6500 7844 6556
rect 7780 6496 7844 6500
rect 7860 6556 7924 6560
rect 7860 6500 7864 6556
rect 7864 6500 7920 6556
rect 7920 6500 7924 6556
rect 7860 6496 7924 6500
rect 7940 6556 8004 6560
rect 7940 6500 7944 6556
rect 7944 6500 8000 6556
rect 8000 6500 8004 6556
rect 7940 6496 8004 6500
rect 13620 6556 13684 6560
rect 13620 6500 13624 6556
rect 13624 6500 13680 6556
rect 13680 6500 13684 6556
rect 13620 6496 13684 6500
rect 13700 6556 13764 6560
rect 13700 6500 13704 6556
rect 13704 6500 13760 6556
rect 13760 6500 13764 6556
rect 13700 6496 13764 6500
rect 13780 6556 13844 6560
rect 13780 6500 13784 6556
rect 13784 6500 13840 6556
rect 13840 6500 13844 6556
rect 13780 6496 13844 6500
rect 13860 6556 13924 6560
rect 13860 6500 13864 6556
rect 13864 6500 13920 6556
rect 13920 6500 13924 6556
rect 13860 6496 13924 6500
rect 13940 6556 14004 6560
rect 13940 6500 13944 6556
rect 13944 6500 14000 6556
rect 14000 6500 14004 6556
rect 13940 6496 14004 6500
<< metal4 >>
rect 6872 13646 7272 13728
rect 6872 13632 6954 13646
rect 7190 13632 7272 13646
rect 6872 13568 6880 13632
rect 6944 13568 6954 13632
rect 7190 13568 7200 13632
rect 7264 13568 7272 13632
rect 6872 13410 6954 13568
rect 7190 13410 7272 13568
rect 6872 12544 7272 13410
rect 6872 12480 6880 12544
rect 6944 12480 6960 12544
rect 7024 12480 7040 12544
rect 7104 12480 7120 12544
rect 7184 12480 7200 12544
rect 7264 12480 7272 12544
rect 6872 11456 7272 12480
rect 6872 11392 6880 11456
rect 6944 11392 6960 11456
rect 7024 11392 7040 11456
rect 7104 11392 7120 11456
rect 7184 11392 7200 11456
rect 7264 11392 7272 11456
rect 6872 10368 7272 11392
rect 6872 10304 6880 10368
rect 6944 10304 6960 10368
rect 7024 10304 7040 10368
rect 7104 10304 7120 10368
rect 7184 10304 7200 10368
rect 7264 10304 7272 10368
rect 6872 9280 7272 10304
rect 6872 9216 6880 9280
rect 6944 9216 6960 9280
rect 7024 9216 7040 9280
rect 7104 9216 7120 9280
rect 7184 9216 7200 9280
rect 7264 9216 7272 9280
rect 6872 8192 7272 9216
rect 6872 8128 6880 8192
rect 6944 8128 6960 8192
rect 7024 8128 7040 8192
rect 7104 8128 7120 8192
rect 7184 8128 7200 8192
rect 7264 8128 7272 8192
rect 6872 7646 7272 8128
rect 6872 7410 6954 7646
rect 7190 7410 7272 7646
rect 6872 7104 7272 7410
rect 6872 7040 6880 7104
rect 6944 7040 6960 7104
rect 7024 7040 7040 7104
rect 7104 7040 7120 7104
rect 7184 7040 7200 7104
rect 7264 7040 7272 7104
rect 6872 6480 7272 7040
rect 7612 13088 8012 13648
rect 7612 13024 7620 13088
rect 7684 13024 7700 13088
rect 7764 13024 7780 13088
rect 7844 13024 7860 13088
rect 7924 13024 7940 13088
rect 8004 13024 8012 13088
rect 7612 12000 8012 13024
rect 7612 11936 7620 12000
rect 7684 11936 7700 12000
rect 7764 11936 7780 12000
rect 7844 11936 7860 12000
rect 7924 11936 7940 12000
rect 8004 11936 8012 12000
rect 7612 10912 8012 11936
rect 7612 10848 7620 10912
rect 7684 10848 7700 10912
rect 7764 10848 7780 10912
rect 7844 10848 7860 10912
rect 7924 10848 7940 10912
rect 8004 10848 8012 10912
rect 7612 9824 8012 10848
rect 7612 9760 7620 9824
rect 7684 9760 7700 9824
rect 7764 9760 7780 9824
rect 7844 9760 7860 9824
rect 7924 9760 7940 9824
rect 8004 9760 8012 9824
rect 7612 8736 8012 9760
rect 7612 8672 7620 8736
rect 7684 8672 7700 8736
rect 7764 8672 7780 8736
rect 7844 8672 7860 8736
rect 7924 8672 7940 8736
rect 8004 8672 8012 8736
rect 7612 8386 8012 8672
rect 7612 8150 7694 8386
rect 7930 8150 8012 8386
rect 7612 7648 8012 8150
rect 7612 7584 7620 7648
rect 7684 7584 7700 7648
rect 7764 7584 7780 7648
rect 7844 7584 7860 7648
rect 7924 7584 7940 7648
rect 8004 7584 8012 7648
rect 7612 6560 8012 7584
rect 7612 6496 7620 6560
rect 7684 6496 7700 6560
rect 7764 6496 7780 6560
rect 7844 6496 7860 6560
rect 7924 6496 7940 6560
rect 8004 6496 8012 6560
rect 7612 6480 8012 6496
rect 12872 13646 13272 13728
rect 12872 13632 12954 13646
rect 13190 13632 13272 13646
rect 12872 13568 12880 13632
rect 12944 13568 12954 13632
rect 13190 13568 13200 13632
rect 13264 13568 13272 13632
rect 12872 13410 12954 13568
rect 13190 13410 13272 13568
rect 12872 12544 13272 13410
rect 12872 12480 12880 12544
rect 12944 12480 12960 12544
rect 13024 12480 13040 12544
rect 13104 12480 13120 12544
rect 13184 12480 13200 12544
rect 13264 12480 13272 12544
rect 12872 11456 13272 12480
rect 12872 11392 12880 11456
rect 12944 11392 12960 11456
rect 13024 11392 13040 11456
rect 13104 11392 13120 11456
rect 13184 11392 13200 11456
rect 13264 11392 13272 11456
rect 12872 10368 13272 11392
rect 12872 10304 12880 10368
rect 12944 10304 12960 10368
rect 13024 10304 13040 10368
rect 13104 10304 13120 10368
rect 13184 10304 13200 10368
rect 13264 10304 13272 10368
rect 12872 9280 13272 10304
rect 12872 9216 12880 9280
rect 12944 9216 12960 9280
rect 13024 9216 13040 9280
rect 13104 9216 13120 9280
rect 13184 9216 13200 9280
rect 13264 9216 13272 9280
rect 12872 8192 13272 9216
rect 12872 8128 12880 8192
rect 12944 8128 12960 8192
rect 13024 8128 13040 8192
rect 13104 8128 13120 8192
rect 13184 8128 13200 8192
rect 13264 8128 13272 8192
rect 12872 7646 13272 8128
rect 12872 7410 12954 7646
rect 13190 7410 13272 7646
rect 12872 7104 13272 7410
rect 12872 7040 12880 7104
rect 12944 7040 12960 7104
rect 13024 7040 13040 7104
rect 13104 7040 13120 7104
rect 13184 7040 13200 7104
rect 13264 7040 13272 7104
rect 12872 6480 13272 7040
rect 13612 13088 14012 13648
rect 13612 13024 13620 13088
rect 13684 13024 13700 13088
rect 13764 13024 13780 13088
rect 13844 13024 13860 13088
rect 13924 13024 13940 13088
rect 14004 13024 14012 13088
rect 13612 12000 14012 13024
rect 13612 11936 13620 12000
rect 13684 11936 13700 12000
rect 13764 11936 13780 12000
rect 13844 11936 13860 12000
rect 13924 11936 13940 12000
rect 14004 11936 14012 12000
rect 13612 10912 14012 11936
rect 13612 10848 13620 10912
rect 13684 10848 13700 10912
rect 13764 10848 13780 10912
rect 13844 10848 13860 10912
rect 13924 10848 13940 10912
rect 14004 10848 14012 10912
rect 13612 9824 14012 10848
rect 13612 9760 13620 9824
rect 13684 9760 13700 9824
rect 13764 9760 13780 9824
rect 13844 9760 13860 9824
rect 13924 9760 13940 9824
rect 14004 9760 14012 9824
rect 13612 8736 14012 9760
rect 13612 8672 13620 8736
rect 13684 8672 13700 8736
rect 13764 8672 13780 8736
rect 13844 8672 13860 8736
rect 13924 8672 13940 8736
rect 14004 8672 14012 8736
rect 13612 8386 14012 8672
rect 13612 8150 13694 8386
rect 13930 8150 14012 8386
rect 13612 7648 14012 8150
rect 13612 7584 13620 7648
rect 13684 7584 13700 7648
rect 13764 7584 13780 7648
rect 13844 7584 13860 7648
rect 13924 7584 13940 7648
rect 14004 7584 14012 7648
rect 13612 6560 14012 7584
rect 13612 6496 13620 6560
rect 13684 6496 13700 6560
rect 13764 6496 13780 6560
rect 13844 6496 13860 6560
rect 13924 6496 13940 6560
rect 14004 6496 14012 6560
rect 13612 6480 14012 6496
<< via4 >>
rect 6954 13632 7190 13646
rect 6954 13568 6960 13632
rect 6960 13568 7024 13632
rect 7024 13568 7040 13632
rect 7040 13568 7104 13632
rect 7104 13568 7120 13632
rect 7120 13568 7184 13632
rect 7184 13568 7190 13632
rect 6954 13410 7190 13568
rect 6954 7410 7190 7646
rect 7694 8150 7930 8386
rect 12954 13632 13190 13646
rect 12954 13568 12960 13632
rect 12960 13568 13024 13632
rect 13024 13568 13040 13632
rect 13040 13568 13104 13632
rect 13104 13568 13120 13632
rect 13120 13568 13184 13632
rect 13184 13568 13190 13632
rect 12954 13410 13190 13568
rect 12954 7410 13190 7646
rect 13694 8150 13930 8386
<< metal5 >>
rect 6024 13646 14032 13728
rect 6024 13410 6954 13646
rect 7190 13410 12954 13646
rect 13190 13410 14032 13646
rect 6024 13328 14032 13410
rect 6024 8386 14032 8468
rect 6024 8150 7694 8386
rect 7930 8150 13694 8386
rect 13930 8150 14032 8386
rect 6024 8068 14032 8150
rect 6024 7646 14032 7728
rect 6024 7410 6954 7646
rect 7190 7410 12954 7646
rect 13190 7410 14032 7646
rect 6024 7328 14032 7410
use sky130_fd_sc_hd__inv_2  _1_
timestamp 0
transform 1 0 7360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2_
timestamp 0
transform 1 0 6716 0 1 9792
box -38 -48 1970 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 8556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 10948 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 11316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_81
timestamp 0
transform 1 0 13524 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 11132 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 12420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_81
timestamp 0
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 8556 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 9844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 10948 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 13156 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 11132 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 12420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_81
timestamp 0
transform 1 0 13524 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 6348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 8556 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 9844 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 10948 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 12052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 13156 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_11
timestamp 0
transform 1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_17
timestamp 0
transform 1 0 7636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_29
timestamp 0
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_41
timestamp 0
transform 1 0 9844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 0
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 12420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_81
timestamp 0
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_6
timestamp 0
transform 1 0 6624 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 9844 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 10948 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 12052 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 13156 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 0
transform 1 0 6624 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_18
timestamp 0
transform 1 0 7728 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_30
timestamp 0
transform 1 0 8832 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_42
timestamp 0
transform 1 0 9936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 0
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_81
timestamp 0
transform 1 0 13524 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 6348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 8556 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 9844 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 13156 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 11132 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 12420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_81
timestamp 0
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 9844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 10948 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 13156 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 11132 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 12420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_81
timestamp 0
transform 1 0 13524 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 8556 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 9844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_53
timestamp 0
transform 1 0 10948 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_57
timestamp 0
transform 1 0 11316 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_69
timestamp 0
transform 1 0 12420 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_81
timestamp 0
transform 1 0 13524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 6624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 0
transform 1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 13984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 0
transform 1 0 6072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 0
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 0
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 13984 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 0
transform 1 0 6072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 0
transform 1 0 6072 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 13984 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 0
transform 1 0 6072 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 0
transform 1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 13984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 0
transform 1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 13984 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 0
transform 1 0 6072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 0
transform 1 0 6072 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 0
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp 0
transform 1 0 11224 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp 0
transform 1 0 11224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp 0
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_30
timestamp 0
transform 1 0 11224 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_31
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_32
timestamp 0
transform 1 0 11224 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_33
timestamp 0
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_34
timestamp 0
transform 1 0 11224 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_35
timestamp 0
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_36
timestamp 0
transform 1 0 11224 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_37
timestamp 0
transform 1 0 8648 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_38
timestamp 0
transform 1 0 11224 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_39
timestamp 0
transform 1 0 8648 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_40
timestamp 0
transform 1 0 11224 0 1 13056
box -38 -48 130 592
<< labels >>
rlabel metal1 s 10042 13056 10042 13056 4 VGND
rlabel metal1 s 10028 13600 10028 13600 4 VPWR
rlabel metal2 s 7498 9826 7498 9826 4 _0_
rlabel metal3 s 2752 9588 2752 9588 4 en
rlabel metal3 s 3534 10268 3534 10268 4 in
rlabel metal1 s 6992 9894 6992 9894 4 net1
rlabel metal2 s 6762 10268 6762 10268 4 net2
rlabel metal2 s 15226 10115 15226 10115 4 out
flabel metal5 s 6024 8068 14032 8468 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 13612 6480 14012 13648 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7612 6480 8012 13648 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 6024 13328 14032 13728 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 6024 7328 14032 7728 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 12872 6480 13272 13728 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 6872 6480 7272 13728 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 en
port 3 nsew
flabel metal3 s 0 10208 800 10328 0 FreeSans 600 0 0 0 in
port 4 nsew
flabel metal3 s 19200 10208 20000 10328 0 FreeSans 600 0 0 0 out
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
